/************************************************************************
	
	fx3StateMachine.v
	FX3 State-Machine module
	
	Domesday Duplicator - LaserDisc RF sampler
	SPDX-FileCopyrightText: 2018-2025 Simon Inns
	SPDX-License-Identifier: GPL-3.0-or-later
	
************************************************************************/

module fx3StateMachine (
	input nReset,
	input fx3_clock,
	input readData,
	
	output fx3isReading
);

// State machine logic ---------------------------------------------------

// State machine state definitions (4-bit 0-15)
reg [3:0]sm_currentState;
reg [3:0]sm_nextState;

parameter [3:0] state_waitForRequest	= 4'd01;
parameter [3:0] state_sendPacket			= 4'd02;

// Set state to state_idle on reset - or assign the next state
always @(posedge fx3_clock, negedge nReset) begin
	if(!nReset) begin 
		sm_currentState <= state_waitForRequest;
	end else begin
		sm_currentState <= sm_nextState;
	end	
end

// Ensure that the readData signal is only read
// on the FX3 clock edge
reg readData_flag;

always @(posedge fx3_clock, negedge nReset) begin
	if(!nReset) begin 
		readData_flag <= 1'b0;
	end else begin
		readData_flag <= readData;
	end	
end

// Counter for the sendPacket state
// Here we should send 8192 words to the FX3
reg [15:0] wordCounter;

always @(posedge fx3_clock, negedge nReset) begin
	if (!nReset) begin
		wordCounter = 16'd0;
	end else begin
		if (sm_currentState == state_sendPacket) begin
			wordCounter = wordCounter + 16'd1;
		end else begin
			wordCounter = 16'd0;
		end
	end
end

// Generate fx3isReading flag
assign fx3isReading = (sm_currentState == state_sendPacket) ? 1'b1 : 1'b0;

// State machine transition logic
always @(*)begin
	sm_nextState = sm_currentState;
	
	case(sm_currentState)
		
		// state_waitForRequest (waits for the FX3 to request a packet)
		state_waitForRequest:begin
			// Is the GPIF reading data?
			if (readData_flag == 1'b1 && wordCounter == 16'd0) begin
				sm_nextState = state_sendPacket;
			end else begin
				// GPIF not ready... wait
				sm_nextState = state_waitForRequest;
			end
		end
		
		// state_sendPacket (sends a packet of 8192 words to the FX3)
		state_sendPacket:begin
			if (wordCounter == 16'd8191) begin
				// Packet send, go back to waiting
				sm_nextState = state_waitForRequest;
			end else begin
				// Continue sending packet
				sm_nextState = state_sendPacket;
			end
		end
		
	endcase
end


endmodule